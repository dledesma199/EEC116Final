magic
tech scmos
timestamp 1702318452
<< ntransistor >>
rect -88 -43 -86 -38
rect -62 -43 -60 -38
rect -35 -43 -33 -38
rect -6 -43 -4 -38
rect 21 -43 23 -38
rect 51 -43 53 -38
rect 81 -43 83 -38
rect 112 -43 114 -38
rect 144 -43 146 -38
rect 176 -43 178 -38
rect 205 -43 207 -38
rect 236 -43 238 -38
rect 270 -43 272 -38
<< ptransistor >>
rect -88 0 -86 5
rect -62 0 -60 5
rect -35 0 -33 5
rect -5 0 -3 5
rect 21 0 23 5
rect 51 0 53 5
rect 81 0 83 5
rect 112 0 114 5
rect 144 0 146 5
rect 176 0 178 5
rect 205 0 207 5
rect 236 0 238 5
rect 270 0 272 5
<< ndiffusion >>
rect -91 -43 -88 -38
rect -86 -43 -81 -38
rect -66 -43 -62 -38
rect -60 -43 -55 -38
rect -39 -43 -35 -38
rect -33 -43 -28 -38
rect -10 -43 -6 -38
rect -4 -43 0 -38
rect 15 -43 21 -38
rect 23 -43 29 -38
rect 45 -43 51 -38
rect 53 -43 59 -38
rect 76 -43 81 -38
rect 83 -43 89 -38
rect 107 -43 112 -38
rect 114 -43 120 -38
rect 138 -43 144 -38
rect 146 -43 152 -38
rect 169 -43 176 -38
rect 178 -43 183 -38
rect 199 -43 205 -38
rect 207 -43 214 -38
rect 230 -43 236 -38
rect 238 -43 244 -38
rect 263 -43 270 -38
rect 272 -43 277 -38
<< pdiffusion >>
rect -91 0 -88 5
rect -86 0 -81 5
rect -65 0 -62 5
rect -60 0 -55 5
rect -39 0 -35 5
rect -33 0 -28 5
rect -10 0 -5 5
rect -3 0 0 5
rect 15 0 21 5
rect 23 0 29 5
rect 45 0 51 5
rect 53 0 59 5
rect 75 0 81 5
rect 83 0 89 5
rect 107 0 112 5
rect 114 0 120 5
rect 138 0 144 5
rect 146 0 152 5
rect 169 0 176 5
rect 178 0 183 5
rect 199 0 205 5
rect 207 0 214 5
rect 230 0 236 5
rect 238 0 244 5
rect 263 0 270 5
rect 272 0 277 5
<< ndcontact >>
rect -96 -43 -91 -38
rect -81 -43 -76 -38
rect -71 -43 -66 -38
rect -55 -43 -50 -38
rect -44 -43 -39 -38
rect -28 -43 -23 -38
rect -15 -43 -10 -38
rect 0 -43 5 -38
rect 10 -43 15 -38
rect 29 -43 34 -38
rect 40 -43 45 -38
rect 59 -43 64 -38
rect 71 -43 76 -38
rect 89 -43 94 -38
rect 102 -43 107 -38
rect 120 -43 125 -38
rect 133 -43 138 -38
rect 152 -43 157 -38
rect 164 -43 169 -38
rect 183 -43 188 -38
rect 194 -43 199 -38
rect 214 -43 219 -38
rect 225 -43 230 -38
rect 244 -43 249 -38
rect 258 -43 263 -38
rect 277 -43 282 -38
<< pdcontact >>
rect -96 0 -91 5
rect -81 0 -76 5
rect -70 0 -65 5
rect -55 0 -50 5
rect -44 0 -39 5
rect -28 0 -23 5
rect -15 0 -10 5
rect 0 0 5 5
rect 10 0 15 5
rect 29 0 34 5
rect 40 0 45 5
rect 59 0 64 5
rect 70 0 75 5
rect 89 0 94 5
rect 102 0 107 5
rect 120 0 125 5
rect 133 0 138 5
rect 152 0 157 5
rect 164 0 169 5
rect 183 0 188 5
rect 194 0 199 5
rect 214 0 219 5
rect 225 0 230 5
rect 244 0 249 5
rect 258 0 263 5
rect 277 0 282 5
<< polysilicon >>
rect -88 5 -86 10
rect -62 5 -60 9
rect -35 5 -33 21
rect -5 5 -3 19
rect 21 5 23 19
rect 51 5 53 19
rect 81 5 83 22
rect 112 5 114 19
rect 144 5 146 19
rect 176 5 178 9
rect 205 5 207 9
rect 236 5 238 9
rect 270 5 272 9
rect -88 -13 -86 0
rect -62 -10 -60 0
rect -35 -3 -33 0
rect -5 -3 -3 0
rect -88 -38 -86 -18
rect -62 -38 -60 -14
rect 21 -19 23 0
rect 51 -8 53 0
rect -35 -38 -33 -34
rect -6 -38 -4 -35
rect 21 -38 23 -23
rect 51 -38 53 -12
rect 81 -28 83 0
rect 112 -3 114 0
rect 144 -3 146 0
rect 176 -16 178 0
rect 205 -16 207 0
rect 236 -16 238 0
rect 270 -15 272 0
rect 81 -38 83 -32
rect 112 -38 114 -33
rect 144 -38 146 -33
rect 176 -38 178 -20
rect 205 -38 207 -20
rect 236 -38 238 -20
rect 270 -38 272 -19
rect -88 -47 -86 -43
rect -62 -47 -60 -43
rect -35 -60 -33 -43
rect -6 -60 -4 -43
rect 21 -48 23 -43
rect 51 -48 53 -43
rect 81 -47 83 -43
rect 112 -57 114 -43
rect 144 -57 146 -43
rect 176 -47 178 -43
rect 205 -47 207 -43
rect 236 -47 238 -43
rect 270 -47 272 -43
<< polycontact >>
rect -37 21 -33 25
rect -6 19 -2 23
rect 111 19 115 23
rect 143 19 147 23
rect -63 -14 -59 -10
rect 50 -12 54 -8
rect 20 -23 24 -19
rect 175 -20 179 -16
rect 204 -20 208 -16
rect 235 -20 239 -16
rect 269 -19 273 -15
rect 80 -32 84 -28
rect -36 -64 -32 -60
rect -7 -64 -3 -60
rect 111 -61 115 -57
rect 143 -61 147 -57
<< metal1 >>
rect -96 47 -50 52
rect -45 47 -37 52
rect -32 47 140 52
rect 145 47 282 52
rect -96 35 -75 40
rect -70 35 282 40
rect -37 25 -33 26
rect -6 23 -2 35
rect 111 23 115 35
rect 140 23 144 27
rect 140 19 143 23
rect -96 8 282 16
rect -96 5 -91 8
rect -70 5 -65 8
rect 10 5 15 8
rect 40 5 45 8
rect 70 5 75 8
rect 164 5 169 8
rect 194 5 199 8
rect 225 5 230 8
rect 258 5 263 8
rect -81 -10 -76 0
rect -81 -14 -63 -10
rect -55 -13 -50 0
rect -81 -23 -76 -14
rect -81 -27 -73 -23
rect -114 -36 -109 -31
rect -81 -38 -76 -27
rect -55 -38 -50 -18
rect -44 -38 -39 0
rect -28 -5 -23 0
rect -15 -5 -10 0
rect -28 -8 -10 -5
rect -28 -18 -23 -8
rect -28 -38 -23 -23
rect -15 -38 -10 -8
rect 0 -5 5 0
rect 0 -38 5 -10
rect 29 -8 34 0
rect 59 -7 64 0
rect 29 -12 50 -8
rect 13 -23 20 -19
rect 29 -27 34 -12
rect 29 -38 34 -32
rect 59 -38 64 -12
rect 89 -13 94 0
rect 102 -13 107 0
rect 89 -19 107 -13
rect 73 -32 80 -28
rect 89 -38 94 -19
rect 102 -38 107 -19
rect 120 -15 125 0
rect 133 -15 138 0
rect 120 -21 138 -15
rect 120 -26 125 -21
rect 120 -38 125 -31
rect 133 -38 138 -21
rect 152 -9 157 0
rect 152 -38 157 -14
rect 183 -16 188 0
rect 214 -8 219 0
rect 166 -21 175 -16
rect 183 -20 204 -16
rect 166 -26 171 -21
rect 183 -27 188 -20
rect 183 -38 188 -32
rect 214 -38 219 -13
rect 244 -15 249 0
rect 226 -20 235 -16
rect 244 -18 269 -15
rect 244 -19 256 -18
rect 226 -27 230 -20
rect 244 -38 249 -19
rect 261 -19 269 -18
rect 277 -38 282 0
rect -96 -46 -91 -43
rect -71 -46 -66 -43
rect 10 -46 15 -43
rect 40 -46 45 -43
rect 71 -46 76 -43
rect 164 -46 169 -43
rect 194 -46 199 -43
rect 225 -46 230 -43
rect 258 -46 263 -43
rect -96 -54 283 -46
rect -36 -73 -32 -64
rect -8 -64 -7 -61
rect 107 -61 111 -59
rect 107 -64 115 -61
rect -8 -65 -4 -64
rect 143 -73 147 -61
rect -96 -78 -75 -73
rect -70 -78 282 -73
rect -96 -89 -50 -84
rect -45 -89 -10 -84
rect -5 -89 107 -84
rect 112 -89 282 -84
<< m2contact >>
rect -50 47 -45 52
rect -37 47 -32 52
rect 140 47 145 52
rect -75 35 -70 40
rect -37 26 -32 31
rect 140 27 145 32
rect -55 -18 -50 -13
rect -73 -28 -68 -23
rect -28 -23 -23 -18
rect 0 -10 5 -5
rect 59 -12 64 -7
rect 8 -23 13 -18
rect 29 -32 34 -27
rect 68 -32 73 -27
rect 120 -31 125 -26
rect 152 -14 157 -9
rect 214 -13 219 -8
rect 166 -31 171 -26
rect 183 -32 188 -27
rect 226 -32 231 -27
rect 256 -23 261 -18
rect -10 -70 -5 -65
rect 107 -69 112 -64
rect -75 -78 -70 -73
rect -50 -89 -45 -84
rect -10 -89 -5 -84
rect 107 -89 112 -84
<< pm12contact >>
rect -91 -18 -86 -13
<< metal2 >>
rect -75 -13 -70 35
rect -101 -18 -91 -13
rect -73 -23 -70 -13
rect -73 -32 -70 -28
rect -75 -73 -70 -32
rect -50 -84 -45 47
rect -37 31 -33 47
rect 140 32 145 47
rect 6 20 69 25
rect 6 -5 11 20
rect 5 -10 11 -5
rect 64 -12 69 20
rect 157 -13 214 -9
rect -23 -23 8 -18
rect 34 -32 68 -27
rect 125 -31 166 -26
rect 188 -32 226 -27
rect 256 -28 293 -23
rect -9 -84 -5 -70
rect 107 -84 112 -69
<< m123contact >>
rect -106 -18 -101 -13
rect -109 -36 -104 -31
rect -39 -22 -34 -17
<< metal3 >>
rect -111 -18 -106 -13
rect -109 -56 -104 -36
rect -39 -56 -34 -22
rect -109 -61 -34 -56
<< m345contact >>
rect -116 -18 -111 -13
<< metal5 >>
rect -126 -18 -116 -13
<< labels >>
rlabel metal1 -53 -24 -53 -24 1 clock_buf
rlabel metal1 -79 -15 -79 -15 1 clock_buf_bar
rlabel metal1 255 -18 255 -18 1 Q
rlabel metal1 279 -16 279 -16 7 Q_NOT
rlabel metal1 -88 11 -88 11 1 Vdd
rlabel metal1 -88 -52 -88 -52 1 Gnd
rlabel metal1 -112 -33 -112 -33 3 D
rlabel metal5 -125 -15 -125 -15 3 CLK
<< end >>
