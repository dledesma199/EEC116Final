magic
tech scmos
timestamp 1702537836
<< metal1 >>
rect -21 1521 0 1529
rect 16 1512 21 1521
rect 66 1496 69 1500
rect 7 1474 10 1478
rect 968 1474 976 1478
rect 421 1464 427 1468
rect 16 1439 21 1447
rect -21 1431 0 1439
rect 426 1415 862 1416
rect 431 1411 862 1415
rect -20 1392 0 1400
rect 16 1383 21 1392
rect 61 1367 69 1371
rect 2 1345 10 1349
rect 968 1345 976 1349
rect 16 1310 21 1318
rect -20 1302 0 1310
rect 426 1286 862 1289
rect 431 1284 862 1286
rect -20 1263 0 1271
rect 16 1254 21 1263
rect 61 1238 69 1242
rect 2 1216 10 1220
rect 968 1217 976 1221
rect 16 1181 21 1189
rect -20 1173 0 1181
rect 431 1152 862 1157
rect -20 1134 0 1142
rect 16 1125 21 1134
rect 61 1109 69 1113
rect 2 1087 10 1091
rect 968 1088 976 1092
rect 16 1052 21 1060
rect -20 1044 0 1052
rect 426 1028 862 1029
rect 431 1024 862 1028
rect -20 1005 0 1013
rect 16 996 21 1005
rect 61 980 69 984
rect 2 958 10 962
rect 968 956 976 960
rect 16 923 21 931
rect -20 915 0 923
rect 426 899 862 900
rect 431 895 862 899
rect -20 876 0 884
rect 16 867 21 876
rect 61 851 69 855
rect 2 829 10 833
rect 968 826 976 830
rect 16 794 21 802
rect -20 786 0 794
rect 426 770 862 771
rect 431 766 862 770
rect -20 747 0 755
rect 16 738 21 747
rect 61 722 69 726
rect 2 700 10 704
rect 968 701 976 705
rect 16 665 21 673
rect -20 657 0 665
rect 426 641 862 642
rect 431 637 862 641
rect -20 618 0 626
rect 16 609 21 618
rect 61 593 69 597
rect 2 571 10 575
rect 968 566 976 570
rect 16 536 21 544
rect -20 528 0 536
rect 426 512 862 513
rect 431 508 862 512
rect -20 489 0 497
rect 16 480 21 489
rect 61 464 69 468
rect 2 442 10 446
rect 968 435 976 439
rect 16 407 21 415
rect -20 399 0 407
rect 426 383 862 384
rect 431 379 862 383
rect -20 360 0 368
rect 16 351 21 360
rect 61 335 69 339
rect 2 313 10 317
rect 968 309 976 313
rect 16 278 21 286
rect -20 270 0 278
rect 426 254 862 255
rect 431 250 862 254
rect -20 231 0 239
rect 16 222 21 231
rect 61 206 69 210
rect 2 184 10 188
rect 968 178 976 182
rect 16 149 21 157
rect -20 141 0 149
rect 426 125 862 126
rect 431 121 862 125
rect -20 102 0 110
rect 16 93 21 102
rect 66 77 69 81
rect 7 55 10 59
rect 968 51 976 55
rect 16 20 21 28
rect -20 12 0 20
rect 431 -11 862 -6
rect -22 -36 0 -28
rect 16 -45 21 -36
rect 857 -63 867 -58
rect 968 -84 976 -80
rect 16 -118 21 -110
rect -22 -126 0 -118
<< m2contact >>
rect 61 77 66 82
rect 2 55 7 60
rect 66 -61 71 -56
rect 7 -83 12 -78
rect 7 -126 12 -121
rect 66 -126 71 -121
<< metal2 >>
rect 7 -121 12 -83
rect 66 -121 71 -61
<< m123contact >>
rect 852 1492 857 1497
rect 426 1410 431 1415
rect 862 1411 867 1416
rect 852 1365 857 1370
rect 426 1335 431 1340
rect 426 1281 431 1286
rect 862 1284 867 1289
rect 852 1233 857 1238
rect 426 1206 431 1211
rect 426 1152 431 1157
rect 862 1152 867 1157
rect 852 1105 857 1110
rect 426 1077 431 1082
rect 426 1023 431 1028
rect 862 1024 867 1029
rect 852 976 857 981
rect 426 948 431 953
rect 426 894 431 899
rect 862 895 867 900
rect 852 847 857 852
rect 426 819 431 824
rect 426 765 431 770
rect 862 766 867 771
rect 852 718 857 723
rect 426 690 431 695
rect 426 636 431 641
rect 862 637 867 642
rect 852 589 857 594
rect 426 561 431 566
rect 426 507 431 512
rect 862 508 867 513
rect 852 460 857 465
rect 426 432 431 437
rect 426 378 431 383
rect 862 379 867 384
rect 852 331 857 336
rect 426 303 431 308
rect 426 249 431 254
rect 862 250 867 255
rect 852 202 857 207
rect 426 174 431 179
rect 426 120 431 125
rect 862 121 867 126
rect 852 76 857 81
rect 426 45 431 50
rect 426 -11 431 -6
rect 862 -11 867 -6
rect 426 -93 431 -88
<< metal3 >>
rect 857 1492 867 1497
rect 862 1416 867 1492
rect 426 1340 431 1410
rect 857 1365 867 1370
rect 862 1289 867 1365
rect 426 1211 431 1281
rect 857 1233 867 1238
rect 862 1157 867 1233
rect 426 1082 431 1152
rect 857 1105 867 1110
rect 862 1029 867 1105
rect 426 953 431 1023
rect 857 976 867 981
rect 862 900 867 976
rect 426 824 431 894
rect 857 847 867 852
rect 862 771 867 847
rect 426 695 431 765
rect 857 718 867 723
rect 862 642 867 718
rect 426 641 431 642
rect 426 566 431 636
rect 857 589 867 594
rect 862 513 867 589
rect 426 512 431 513
rect 426 437 431 507
rect 857 460 867 465
rect 862 384 867 460
rect 426 383 431 384
rect 426 308 431 378
rect 857 331 867 336
rect 862 255 867 331
rect 426 254 431 255
rect 426 179 431 249
rect 857 202 867 207
rect 862 126 867 202
rect 426 125 431 126
rect 426 50 431 120
rect 857 76 867 81
rect 862 -6 867 76
rect 426 -88 431 -11
use RCAcomp  RCAcomp_0
array 0 0 1 0 11 129
timestamp 1701901221
transform 1 0 69 0 1 0
box -69 0 899 118
use RCAcomp  RCAcomp_1
timestamp 1701901221
transform 1 0 69 0 1 -138
box -69 0 899 118
<< labels >>
rlabel metal1 -15 1526 -15 1526 1 Vdd
rlabel metal1 -14 1396 -14 1396 1 Vdd
rlabel metal1 -18 1267 -18 1267 3 Vdd
rlabel metal1 -18 1137 -18 1137 3 Vdd
rlabel metal1 -18 1011 -18 1011 3 Vdd
rlabel metal1 -19 882 -19 882 3 Vdd
rlabel metal1 -19 754 -19 754 3 Vdd
rlabel metal1 -19 621 -19 621 3 Vdd
rlabel metal1 -19 492 -19 492 3 Vdd
rlabel metal1 -17 365 -17 365 3 Vdd
rlabel metal1 -18 236 -18 236 3 Vdd
rlabel metal1 -18 106 -18 106 3 Vdd
rlabel metal1 -19 16 -19 16 3 Gnd
rlabel metal1 -17 147 -17 147 3 Gnd
rlabel metal1 -18 274 -18 274 3 Gnd
rlabel metal1 -18 403 -18 403 3 Gnd
rlabel metal1 -18 530 -18 530 3 Gnd
rlabel metal1 -14 659 -14 659 1 Gnd
rlabel metal1 -18 790 -18 790 3 Gnd
rlabel metal1 -16 918 -16 918 3 Gnd
rlabel metal1 -18 1045 -18 1045 3 Gnd
rlabel metal1 -18 1176 -18 1176 3 Gnd
rlabel metal1 -18 1306 -18 1306 3 Gnd
rlabel metal1 -19 1435 -19 1435 3 Gnd
rlabel metal1 423 1467 423 1467 1 Cin0
rlabel metal1 7 1476 7 1476 1 b0
rlabel metal1 66 1497 66 1497 1 a0
rlabel metal1 974 1476 974 1476 7 sum0
rlabel metal1 973 1346 973 1346 7 sum1
rlabel metal1 975 1219 975 1219 7 sum2
rlabel metal1 975 1089 975 1089 7 sum3
rlabel metal1 974 958 974 958 7 sum4
rlabel metal1 974 828 974 828 7 sum5
rlabel metal1 974 703 974 703 7 sum6
rlabel metal1 975 568 975 568 7 sum7
rlabel metal1 975 436 975 436 7 sum8
rlabel metal1 974 311 974 311 7 sum9
rlabel metal1 974 181 974 181 7 sum10
rlabel metal1 975 54 975 54 7 sum11
rlabel metal1 62 1369 62 1369 1 a1
rlabel metal1 4 1347 4 1347 1 b1
rlabel metal1 62 1239 62 1239 1 a2
rlabel metal1 3 1218 3 1218 1 b2
rlabel metal1 62 1111 62 1111 1 a3
rlabel metal1 3 1089 3 1089 1 b3
rlabel metal1 62 982 62 982 1 a4
rlabel metal1 3 960 3 960 1 b4
rlabel metal1 62 853 62 853 1 a5
rlabel metal1 3 831 3 831 1 b5
rlabel metal1 62 724 62 724 1 a6
rlabel metal1 3 702 3 702 1 b6
rlabel metal1 62 595 62 595 1 a7
rlabel metal1 3 573 3 573 1 b7
rlabel metal1 62 466 62 466 1 a8
rlabel metal1 3 444 3 444 1 b8
rlabel metal1 62 337 62 337 1 a9
rlabel metal1 3 315 3 315 1 b9
rlabel metal1 62 208 62 208 1 a10
rlabel metal1 3 186 3 186 1 b10
rlabel m2contact 62 79 62 79 1 a11
rlabel m2contact 3 57 3 57 1 b11
rlabel metal1 974 -82 974 -82 7 sum12
rlabel metal1 865 -61 865 -61 1 Cout12
rlabel metal1 -21 -122 -21 -122 3 Gnd
rlabel metal1 -20 -31 -20 -31 3 Vdd
<< end >>
