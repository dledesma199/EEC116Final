magic
tech scmos
timestamp 1702320260
<< m3contact >>
rect 429 1678 434 1683
rect 429 1531 434 1536
rect 429 1384 434 1389
rect 429 1237 434 1242
rect 429 1090 434 1095
rect 429 943 434 948
rect 429 796 434 801
rect 429 649 434 654
rect 429 502 434 507
rect 429 355 434 360
rect 429 208 434 213
rect 429 61 434 66
<< metal3 >>
rect 434 1678 533 1683
rect 434 1531 524 1536
rect 434 1384 515 1389
rect 434 1237 506 1242
rect 434 1090 497 1095
rect 434 943 488 948
rect 434 796 479 801
rect 434 649 470 654
rect 434 502 461 507
rect 434 355 452 360
rect 434 208 443 213
rect 429 0 434 61
rect 438 0 443 208
rect 447 0 452 355
rect 456 0 461 502
rect 465 0 470 649
rect 474 0 479 796
rect 483 0 488 943
rect 492 0 497 1090
rect 501 0 506 1237
rect 510 0 515 1384
rect 519 0 524 1531
rect 528 0 533 1678
use 12bitRegister  12bitRegister_0
timestamp 1702318452
transform 1 0 15 0 1 0
box -15 0 419 1758
<< end >>
