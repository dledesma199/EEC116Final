magic
tech scmos
timestamp 1702508064
<< nwell >>
rect -6 -27 249 22
rect -6 -30 248 -27
<< pwell >>
rect -6 -67 246 -32
<< ntransistor >>
rect 7 -55 9 -49
rect 40 -54 42 -45
rect 51 -54 53 -45
rect 84 -56 86 -38
rect 95 -56 97 -38
rect 106 -56 108 -38
rect 139 -56 141 -38
rect 150 -56 152 -38
rect 161 -56 163 -38
rect 172 -56 174 -38
rect 183 -56 185 -38
rect 194 -56 196 -38
rect 205 -56 207 -38
rect 216 -56 218 -38
rect 227 -56 229 -38
<< ptransistor >>
rect 7 0 9 12
rect 40 -6 42 12
rect 51 -6 53 12
rect 84 -24 86 12
rect 95 -24 97 12
rect 106 -24 108 12
rect 139 -24 141 12
rect 150 -24 152 12
rect 161 -24 163 12
rect 172 -24 174 12
rect 183 -24 185 12
rect 194 -24 196 12
rect 205 -24 207 12
rect 216 -24 218 12
rect 227 -24 229 12
<< ndiffusion >>
rect 33 -49 40 -45
rect 0 -50 7 -49
rect 5 -55 7 -50
rect 9 -54 11 -49
rect 38 -54 40 -49
rect 42 -50 44 -45
rect 49 -50 51 -45
rect 42 -54 51 -50
rect 53 -49 60 -45
rect 53 -54 55 -49
rect 77 -49 84 -38
rect 82 -54 84 -49
rect 9 -55 16 -54
rect 77 -56 84 -54
rect 86 -43 88 -38
rect 93 -43 95 -38
rect 86 -56 95 -43
rect 97 -49 106 -38
rect 97 -54 99 -49
rect 104 -54 106 -49
rect 97 -56 106 -54
rect 108 -43 110 -38
rect 108 -56 115 -43
rect 132 -51 139 -38
rect 137 -56 139 -51
rect 141 -43 143 -38
rect 148 -43 150 -38
rect 141 -56 150 -43
rect 152 -49 161 -38
rect 152 -54 154 -49
rect 159 -54 161 -49
rect 152 -56 161 -54
rect 163 -43 165 -38
rect 170 -43 172 -38
rect 163 -56 172 -43
rect 174 -49 183 -38
rect 174 -54 176 -49
rect 181 -54 183 -49
rect 174 -56 183 -54
rect 185 -43 187 -38
rect 192 -43 194 -38
rect 185 -56 194 -43
rect 196 -49 205 -38
rect 196 -54 198 -49
rect 203 -54 205 -49
rect 196 -56 205 -54
rect 207 -43 209 -38
rect 214 -43 216 -38
rect 207 -56 216 -43
rect 218 -49 227 -38
rect 218 -54 220 -49
rect 225 -54 227 -49
rect 218 -56 227 -54
rect 229 -43 231 -38
rect 229 -56 236 -43
<< pdiffusion >>
rect 5 7 7 12
rect 0 0 7 7
rect 9 5 16 12
rect 9 0 11 5
rect 38 7 40 12
rect 33 -6 40 7
rect 42 -1 51 12
rect 42 -6 44 -1
rect 49 -6 51 -1
rect 53 7 55 12
rect 53 -6 60 7
rect 82 7 84 12
rect 77 -24 84 7
rect 86 -19 95 12
rect 86 -24 88 -19
rect 93 -24 95 -19
rect 97 7 99 12
rect 104 7 106 12
rect 97 -24 106 7
rect 108 -19 115 12
rect 108 -24 110 -19
rect 137 7 139 12
rect 132 -24 139 7
rect 141 -19 150 12
rect 141 -24 143 -19
rect 148 -24 150 -19
rect 152 7 154 12
rect 159 7 161 12
rect 152 -24 161 7
rect 163 -19 172 12
rect 163 -24 165 -19
rect 170 -24 172 -19
rect 174 7 176 12
rect 181 7 183 12
rect 174 -24 183 7
rect 185 -19 194 12
rect 185 -24 187 -19
rect 192 -24 194 -19
rect 196 7 198 12
rect 203 7 205 12
rect 196 -24 205 7
rect 207 -19 216 12
rect 207 -24 209 -19
rect 214 -24 216 -19
rect 218 7 220 12
rect 225 7 227 12
rect 218 -24 227 7
rect 229 -19 236 12
rect 229 -24 231 -19
<< ndcontact >>
rect 0 -55 5 -50
rect 11 -54 16 -49
rect 33 -54 38 -49
rect 44 -50 49 -45
rect 55 -54 60 -49
rect 77 -54 82 -49
rect 88 -43 93 -38
rect 99 -54 104 -49
rect 110 -43 115 -38
rect 132 -56 137 -51
rect 143 -43 148 -38
rect 154 -54 159 -49
rect 165 -43 170 -38
rect 176 -54 181 -49
rect 187 -43 192 -38
rect 198 -54 203 -49
rect 209 -43 214 -38
rect 220 -54 225 -49
rect 231 -43 236 -38
<< pdcontact >>
rect 0 7 5 12
rect 11 0 16 5
rect 33 7 38 12
rect 44 -6 49 -1
rect 55 7 60 12
rect 77 7 82 12
rect 88 -24 93 -19
rect 99 7 104 12
rect 110 -24 115 -19
rect 132 7 137 12
rect 143 -24 148 -19
rect 154 7 159 12
rect 165 -24 170 -19
rect 176 7 181 12
rect 187 -24 192 -19
rect 198 7 203 12
rect 209 -24 214 -19
rect 220 7 225 12
rect 231 -24 236 -19
<< psubstratepcontact >>
rect 20 -64 25 -59
rect 64 -64 69 -59
rect 121 -64 126 -59
<< nsubstratencontact >>
rect 22 13 27 18
rect 66 13 71 18
rect 120 14 125 19
<< polysilicon >>
rect 7 12 9 15
rect 40 12 42 23
rect 51 12 53 23
rect 84 12 86 23
rect 95 12 97 23
rect 106 12 108 23
rect 139 12 141 23
rect 150 12 152 23
rect 161 12 163 23
rect 172 12 174 23
rect 183 12 185 23
rect 194 12 196 23
rect 205 12 207 23
rect 216 12 218 23
rect 227 12 229 23
rect 7 -16 9 0
rect 40 -15 42 -6
rect 8 -21 9 -16
rect 41 -20 42 -15
rect 7 -49 9 -21
rect 40 -45 42 -20
rect 51 -45 53 -6
rect 84 -26 86 -24
rect 85 -31 86 -26
rect 84 -38 86 -31
rect 95 -38 97 -24
rect 106 -38 108 -24
rect 139 -28 141 -24
rect 140 -33 141 -28
rect 139 -38 141 -33
rect 150 -38 152 -24
rect 161 -38 163 -24
rect 172 -38 174 -24
rect 183 -38 185 -24
rect 194 -38 196 -24
rect 205 -38 207 -24
rect 216 -38 218 -24
rect 227 -38 229 -24
rect 7 -59 9 -55
rect 40 -57 42 -54
rect 51 -57 53 -54
rect 84 -59 86 -56
rect 95 -59 97 -56
rect 106 -59 108 -56
rect 139 -59 141 -56
rect 150 -59 152 -56
rect 161 -59 163 -56
rect 172 -60 174 -56
rect 183 -60 185 -56
rect 194 -59 196 -56
rect 205 -59 207 -56
rect 216 -59 218 -56
rect 227 -59 229 -56
<< polycontact >>
rect 3 -21 8 -16
rect 36 -20 41 -15
rect 80 -31 85 -26
rect 135 -33 140 -28
<< metal1 >>
rect 0 19 236 20
rect 0 18 120 19
rect 0 13 22 18
rect 27 13 66 18
rect 71 14 120 18
rect 125 14 236 19
rect 71 13 236 14
rect 0 12 236 13
rect 11 -15 16 0
rect -11 -21 3 -16
rect 11 -20 36 -15
rect 11 -49 16 -20
rect 44 -26 49 -6
rect 44 -31 80 -26
rect 88 -27 93 -24
rect 110 -27 115 -24
rect 88 -28 115 -27
rect 143 -28 148 -24
rect 165 -28 170 -24
rect 187 -28 192 -24
rect 209 -28 214 -24
rect 231 -28 236 -24
rect 44 -45 49 -31
rect 88 -32 135 -28
rect 88 -38 93 -32
rect 110 -33 135 -32
rect 143 -33 240 -28
rect 110 -38 115 -33
rect 143 -38 148 -33
rect 165 -38 170 -33
rect 187 -38 192 -33
rect 209 -38 214 -33
rect 231 -38 236 -33
rect 0 -58 5 -55
rect 33 -58 38 -54
rect 55 -58 60 -54
rect 77 -58 82 -54
rect 99 -58 104 -54
rect 132 -58 137 -56
rect 154 -58 159 -54
rect 176 -58 181 -54
rect 198 -58 203 -54
rect 220 -58 225 -54
rect 0 -59 236 -58
rect 0 -64 20 -59
rect 25 -64 64 -59
rect 69 -64 121 -59
rect 126 -64 236 -59
rect 0 -66 236 -64
<< pm12contact >>
rect 39 23 44 28
rect 50 23 55 28
rect 82 23 87 28
rect 94 23 99 28
rect 104 23 109 28
rect 138 23 143 28
rect 149 23 154 28
rect 160 23 165 28
rect 170 23 175 28
rect 182 23 187 28
rect 193 23 198 28
rect 204 23 209 28
rect 214 23 219 28
rect 226 23 231 28
<< metal2 >>
rect 44 23 50 28
rect 87 23 94 28
rect 99 23 104 28
rect 143 23 149 28
rect 154 23 160 28
rect 165 23 170 28
rect 175 23 182 28
rect 187 23 193 28
rect 198 23 204 28
rect 209 23 214 28
rect 219 23 226 28
<< end >>
