magic
tech scmos
timestamp 1702571561
<< metal1 >>
rect 962 3417 1121 3425
rect 963 3355 1122 3363
rect 962 3270 1121 3278
rect 963 3208 1122 3216
rect 962 3123 1121 3131
rect 963 3061 1122 3069
rect 962 2976 1121 2984
rect 963 2914 1122 2922
rect 962 2829 1121 2837
rect 963 2767 1122 2775
rect 962 2682 1121 2690
rect 963 2620 1122 2628
rect 962 2535 1121 2543
rect 963 2473 1122 2481
rect 962 2388 1121 2396
rect 963 2326 1122 2334
rect 962 2241 1121 2249
rect 963 2179 1122 2187
rect 962 2094 1121 2102
rect 963 2032 1122 2040
rect 962 1947 1121 1955
rect 963 1885 1122 1893
rect 962 1800 1121 1808
rect 963 1738 1122 1746
rect 1049 1666 1132 1674
rect 1049 1576 1132 1584
rect 1048 1537 1132 1545
rect 1048 1447 1132 1455
rect 1048 1408 1132 1416
rect 1048 1318 1132 1326
rect 1048 1279 1132 1287
rect 1048 1189 1132 1197
rect 1048 1150 1132 1158
rect 1048 1060 1132 1068
rect 1048 1021 1132 1029
rect 1048 931 1132 939
rect 1048 892 1132 900
rect 1048 802 1132 810
rect 1048 763 1132 771
rect 1048 673 1132 681
rect 1048 634 1132 642
rect 1048 544 1132 552
rect 1048 505 1132 513
rect 1048 415 1132 423
rect 1048 376 1132 384
rect 1048 286 1132 294
rect 1048 247 1132 255
rect 1048 157 1132 165
rect 1050 109 1134 117
rect 42 61 61 66
rect 1124 61 1133 66
rect 1050 19 1134 27
<< m2contact >>
rect 1098 3373 1103 3378
rect 1098 3226 1103 3231
rect 1098 3079 1103 3084
rect 1098 2932 1103 2937
rect 1098 2785 1103 2790
rect 1098 2638 1103 2643
rect 1098 2491 1103 2496
rect 1098 2344 1103 2349
rect 1098 2197 1103 2202
rect 1098 2050 1103 2055
rect 1098 1903 1103 1908
rect 1098 1756 1103 1761
rect 1119 61 1124 66
rect 569 -1934 574 -1929
rect 927 -1962 932 -1957
rect 982 -1984 987 -1979
rect 569 -1994 574 -1989
rect 932 -2091 937 -2086
rect 988 -2113 993 -2108
rect 930 -2220 935 -2215
rect 991 -2242 996 -2237
rect 931 -2349 936 -2344
rect 991 -2371 996 -2366
rect 931 -2478 936 -2473
rect 989 -2500 994 -2495
rect 930 -2607 935 -2602
rect 991 -2629 996 -2624
rect 927 -2736 932 -2731
rect 991 -2758 996 -2753
rect 932 -2865 937 -2860
rect 992 -2887 997 -2882
rect 930 -2994 935 -2989
rect 991 -3016 996 -3011
rect 931 -3123 936 -3118
rect 991 -3145 996 -3140
rect 931 -3252 936 -3247
rect 990 -3274 995 -3269
rect 14 -3542 19 -3537
<< metal2 >>
rect 968 3378 973 3386
rect 968 3373 1098 3378
rect 968 3231 973 3239
rect 968 3226 1098 3231
rect 968 3084 973 3092
rect 968 3079 1098 3084
rect 968 2937 973 2945
rect 968 2932 1098 2937
rect 968 2790 973 2798
rect 968 2785 1098 2790
rect 968 2643 973 2651
rect 968 2638 1098 2643
rect 968 2496 973 2504
rect 968 2491 1098 2496
rect 968 2349 973 2357
rect 968 2344 1098 2349
rect 968 2202 973 2210
rect 968 2197 1098 2202
rect 968 2055 973 2063
rect 968 2050 1098 2055
rect 968 1908 973 1916
rect 968 1903 1098 1908
rect 968 1761 973 1769
rect 968 1756 1098 1761
rect 1114 61 1119 66
rect 1868 -660 2139 -655
rect 1868 -669 2031 -664
rect 1868 -736 2022 -731
rect 1868 -745 2130 -740
rect 1868 -758 2121 -753
rect 1868 -767 2013 -762
rect 1868 -834 2004 -829
rect 1868 -843 2112 -838
rect 1868 -856 2103 -851
rect 1868 -865 1995 -860
rect 1868 -932 1986 -927
rect 1868 -941 2094 -936
rect 1868 -954 2085 -949
rect 1868 -963 1977 -958
rect 1868 -1030 1968 -1025
rect 1868 -1039 2076 -1034
rect 1868 -1052 2067 -1047
rect 1868 -1061 1959 -1056
rect 1868 -1128 1950 -1123
rect 1868 -1137 2058 -1132
rect 1868 -1150 2049 -1145
rect 1867 -1159 1941 -1154
rect 1868 -1226 1932 -1221
rect 1868 -1235 2040 -1230
rect 569 -1989 574 -1934
rect 932 -1962 1067 -1957
rect 987 -1984 1076 -1979
rect 934 -2086 1063 -2085
rect 937 -2091 1058 -2086
rect 993 -2113 1085 -2108
rect 935 -2220 1049 -2215
rect 996 -2242 1094 -2237
rect 936 -2349 1040 -2344
rect 996 -2371 1103 -2366
rect 1081 -2430 1205 -2425
rect 1072 -2439 1205 -2434
rect 936 -2478 1031 -2473
rect 989 -2495 1112 -2490
rect 1063 -2506 1205 -2501
rect 1090 -2515 1205 -2510
rect 1099 -2528 1206 -2523
rect 1054 -2537 1205 -2532
rect 935 -2607 1022 -2602
rect 1045 -2604 1205 -2599
rect 1108 -2613 1205 -2608
rect 996 -2641 1001 -2624
rect 1117 -2626 1205 -2621
rect 1036 -2635 1205 -2630
rect 996 -2646 1121 -2641
rect 1027 -2702 1206 -2697
rect 1126 -2711 1205 -2706
rect 1135 -2724 1205 -2719
rect 1018 -2733 1205 -2728
rect 927 -2739 932 -2736
rect 927 -2744 1013 -2739
rect 996 -2758 1130 -2753
rect 1009 -2800 1205 -2795
rect 1144 -2809 1205 -2804
rect 1153 -2822 1205 -2817
rect 1000 -2831 1205 -2826
rect 937 -2865 1004 -2860
rect 997 -2887 1139 -2882
rect 991 -2898 1205 -2893
rect 1162 -2907 1205 -2902
rect 1171 -2920 1205 -2915
rect 982 -2929 1205 -2924
rect 930 -2977 995 -2972
rect 930 -2989 935 -2977
rect 973 -2996 1205 -2991
rect 1180 -3005 1205 -3000
rect 996 -3016 1148 -3011
rect 936 -3123 986 -3118
rect 996 -3145 1157 -3140
rect 936 -3252 977 -3247
rect 995 -3274 1166 -3269
rect 934 -3381 968 -3376
rect 988 -3471 993 -3403
rect 9 -3542 14 -3537
<< m3contact >>
rect 2139 -660 2144 -655
rect 277 -669 282 -664
rect 2031 -669 2036 -664
rect 280 -736 285 -731
rect 2022 -736 2027 -731
rect 2130 -745 2135 -740
rect 2121 -758 2126 -753
rect 275 -767 280 -762
rect 2013 -767 2018 -762
rect 275 -834 280 -829
rect 2004 -834 2009 -829
rect 2112 -843 2117 -838
rect 2103 -856 2108 -851
rect 275 -865 280 -860
rect 1995 -865 2000 -860
rect 275 -932 280 -927
rect 1986 -932 1991 -927
rect 2094 -941 2099 -936
rect 2085 -954 2090 -949
rect 275 -963 280 -958
rect 1977 -963 1982 -958
rect 275 -1030 280 -1025
rect 1968 -1030 1973 -1025
rect 2076 -1039 2081 -1034
rect 2067 -1052 2072 -1047
rect 275 -1061 280 -1056
rect 1959 -1061 1964 -1056
rect 275 -1128 280 -1123
rect 1950 -1128 1955 -1123
rect 2058 -1137 2063 -1132
rect 2049 -1150 2054 -1145
rect 275 -1159 280 -1154
rect 1941 -1159 1946 -1154
rect 275 -1226 280 -1221
rect 1932 -1226 1937 -1221
rect 2040 -1235 2045 -1230
rect 1067 -1962 1072 -1957
rect 1076 -1984 1081 -1979
rect 1058 -2091 1063 -2086
rect 1085 -2113 1090 -2108
rect 1049 -2220 1054 -2215
rect 1094 -2242 1099 -2237
rect 1040 -2349 1045 -2344
rect 1103 -2371 1108 -2366
rect 1076 -2430 1081 -2425
rect 1067 -2439 1072 -2434
rect 1112 -2495 1117 -2490
rect 1058 -2506 1063 -2501
rect 1085 -2515 1090 -2510
rect 1094 -2528 1099 -2523
rect 1049 -2537 1054 -2532
rect 1040 -2604 1045 -2599
rect 1103 -2613 1108 -2608
rect 1112 -2626 1117 -2621
rect 1121 -2646 1126 -2641
rect 1121 -2711 1126 -2706
rect 1130 -2724 1135 -2719
rect 1130 -2758 1135 -2753
rect 1139 -2809 1144 -2804
rect 1148 -2822 1153 -2817
rect 1139 -2887 1144 -2882
rect 1157 -2907 1162 -2902
rect 1166 -2920 1171 -2915
rect 1175 -3005 1180 -3000
rect 1148 -3016 1153 -3011
rect 1157 -3145 1162 -3140
rect 1166 -3274 1171 -3269
rect 988 -3476 993 -3471
<< m123contact >>
rect 37 61 42 66
<< metal3 >>
rect 32 61 37 66
rect 433 -2 438 2
rect 156 -7 438 -2
rect 156 -1221 161 -7
rect 442 -11 447 2
rect 166 -16 447 -11
rect 166 -1154 171 -16
rect 451 -20 456 2
rect 176 -25 456 -20
rect 176 -1123 181 -25
rect 460 -29 465 2
rect 186 -34 465 -29
rect 186 -1056 191 -34
rect 469 -38 474 2
rect 196 -43 474 -38
rect 196 -1025 201 -43
rect 478 -47 483 2
rect 206 -52 483 -47
rect 206 -958 211 -52
rect 487 -56 492 2
rect 216 -61 492 -56
rect 216 -927 221 -61
rect 496 -66 501 2
rect 226 -70 501 -66
rect 226 -860 231 -70
rect 505 -74 510 2
rect 236 -79 510 -74
rect 236 -829 241 -79
rect 514 -83 519 2
rect 246 -88 519 -83
rect 246 -762 251 -88
rect 523 -92 528 2
rect 256 -97 528 -92
rect 256 -731 261 -97
rect 532 -102 537 2
rect 1505 -97 1510 2
rect 1514 -88 1519 2
rect 1523 -79 1528 2
rect 1532 -70 1537 2
rect 1541 -61 1546 2
rect 1550 -52 1555 2
rect 1559 -43 1564 2
rect 1568 -34 1573 2
rect 1577 -25 1582 2
rect 1586 -16 1591 2
rect 1595 -7 1600 2
rect 1604 -3 2036 2
rect 1595 -12 2027 -7
rect 1586 -21 2018 -16
rect 1577 -30 2009 -25
rect 1568 -39 2000 -34
rect 1559 -48 1991 -43
rect 1550 -57 1982 -52
rect 1541 -66 1973 -61
rect 1532 -75 1964 -70
rect 1523 -84 1955 -79
rect 1514 -93 1946 -88
rect 1505 -102 1937 -97
rect 266 -107 537 -102
rect 266 -664 271 -107
rect 266 -669 277 -664
rect 256 -736 280 -731
rect 246 -767 275 -762
rect 236 -834 275 -829
rect 226 -865 275 -860
rect 216 -932 275 -927
rect 206 -963 275 -958
rect 196 -1030 275 -1025
rect 186 -1061 275 -1056
rect 176 -1128 275 -1123
rect 166 -1159 275 -1154
rect 1932 -1221 1937 -102
rect 156 -1226 275 -1221
rect 1932 -1235 1937 -1226
rect 1941 -1154 1946 -93
rect 1941 -1235 1946 -1159
rect 1950 -1123 1955 -84
rect 1950 -1235 1955 -1128
rect 1959 -1056 1964 -75
rect 1959 -1235 1964 -1061
rect 1968 -1025 1973 -66
rect 1968 -1235 1973 -1030
rect 1977 -958 1982 -57
rect 1977 -1235 1982 -963
rect 1986 -927 1991 -48
rect 1986 -1235 1991 -932
rect 1995 -860 2000 -39
rect 1995 -1235 2000 -865
rect 2004 -829 2009 -30
rect 2004 -1235 2009 -834
rect 2013 -762 2018 -21
rect 2013 -1235 2018 -767
rect 2022 -731 2027 -12
rect 2022 -1235 2027 -736
rect 2031 -664 2036 -3
rect 2031 -1235 2036 -669
rect 2040 -1230 2045 2
rect 2049 -1145 2054 2
rect 2058 -1132 2063 2
rect 2067 -1047 2072 2
rect 2076 -1034 2081 3
rect 2085 -949 2090 2
rect 2094 -936 2099 2
rect 2103 -851 2108 2
rect 2112 -838 2117 2
rect 2121 -753 2126 2
rect 2130 -740 2135 2
rect 2139 -655 2144 2
rect 1040 -2344 1045 -1866
rect 1040 -2599 1045 -2349
rect 1040 -3421 1045 -2604
rect 1049 -2215 1054 -1866
rect 1049 -2532 1054 -2220
rect 1049 -3421 1054 -2537
rect 1058 -2086 1063 -1866
rect 1058 -2501 1063 -2091
rect 1058 -3421 1063 -2506
rect 1067 -1957 1072 -1866
rect 1067 -2434 1072 -1962
rect 1067 -3421 1072 -2439
rect 1076 -1979 1081 -1866
rect 1076 -2425 1081 -1984
rect 1076 -3421 1081 -2430
rect 1085 -2108 1090 -1866
rect 1085 -2510 1090 -2113
rect 1085 -3421 1090 -2515
rect 1094 -2237 1099 -1866
rect 1094 -2523 1099 -2242
rect 1094 -3421 1099 -2528
rect 1103 -2366 1108 -1866
rect 1103 -2608 1108 -2371
rect 1103 -3421 1108 -2613
rect 1112 -2490 1117 -1866
rect 1112 -2621 1117 -2495
rect 1112 -3421 1117 -2626
rect 1121 -2641 1126 -1866
rect 1121 -2706 1126 -2646
rect 1121 -3421 1126 -2711
rect 1130 -2719 1135 -1866
rect 1130 -2753 1135 -2724
rect 1130 -3421 1135 -2758
rect 1139 -2804 1144 -1866
rect 1139 -2882 1144 -2809
rect 1139 -3421 1144 -2887
rect 1148 -2817 1153 -1866
rect 1148 -3011 1153 -2822
rect 1148 -3421 1153 -3016
rect 1157 -2902 1162 -1866
rect 1157 -3140 1162 -2907
rect 1157 -3421 1162 -3145
rect 1166 -2915 1171 -1866
rect 1166 -3269 1171 -2920
rect 1166 -3421 1171 -3274
rect 1175 -3000 1180 -1866
rect 1175 -3471 1180 -3005
rect 993 -3476 1180 -3471
<< m234contact >>
rect 1109 61 1114 66
rect 277 -660 282 -655
rect 279 -745 284 -740
rect 275 -758 280 -753
rect 275 -843 280 -838
rect 275 -856 280 -851
rect 275 -941 280 -936
rect 275 -954 280 -949
rect 275 -1039 280 -1034
rect 275 -1052 280 -1047
rect 275 -1137 280 -1132
rect 275 -1150 280 -1145
rect 275 -1235 280 -1230
rect 1031 -2478 1036 -2473
rect 1022 -2607 1027 -2602
rect 1031 -2635 1036 -2630
rect 1022 -2702 1027 -2697
rect 1013 -2733 1018 -2728
rect 1013 -2744 1018 -2739
rect 1004 -2800 1009 -2795
rect 995 -2831 1000 -2826
rect 1004 -2865 1009 -2860
rect 986 -2898 991 -2893
rect 977 -2929 982 -2924
rect 995 -2977 1000 -2972
rect 968 -2996 973 -2991
rect 986 -3123 991 -3118
rect 977 -3252 982 -3247
rect 968 -3381 973 -3376
rect 4 -3542 9 -3537
<< m4contact >>
rect 968 2 973 7
rect 977 2 982 7
rect 986 2 991 7
rect 995 2 1000 7
rect 1004 2 1009 7
rect 1013 2 1018 7
rect 1022 2 1027 7
rect 1031 2 1036 7
rect 1040 2 1045 7
rect 1049 2 1054 7
rect 1058 2 1063 7
rect 1067 2 1072 7
rect 968 -1871 973 -1866
rect 977 -1871 982 -1866
rect 986 -1871 991 -1866
rect 995 -1871 1000 -1866
rect 1004 -1871 1009 -1866
rect 1013 -1871 1018 -1866
rect 1022 -1871 1027 -1866
rect 1031 -1871 1036 -1866
<< metal4 >>
rect 151 -3 973 2
rect 151 -1230 156 -3
rect 977 -7 982 2
rect 161 -12 982 -7
rect 161 -1145 166 -12
rect 986 -16 991 2
rect 171 -21 991 -16
rect 171 -1132 176 -21
rect 995 -25 1000 2
rect 181 -30 1000 -25
rect 181 -1047 186 -30
rect 1004 -34 1009 2
rect 191 -39 1009 -34
rect 191 -1034 196 -39
rect 1013 -43 1018 2
rect 201 -48 1018 -43
rect 201 -949 206 -48
rect 1022 -52 1027 2
rect 211 -57 1027 -52
rect 211 -936 216 -57
rect 1031 -61 1036 2
rect 221 -66 1036 -61
rect 221 -851 226 -66
rect 1040 -70 1045 2
rect 231 -75 1045 -70
rect 231 -838 236 -75
rect 1049 -79 1054 2
rect 241 -84 1054 -79
rect 241 -753 246 -84
rect 1058 -88 1063 2
rect 251 -93 1063 -88
rect 251 -740 256 -93
rect 1067 -97 1072 2
rect 261 -102 1072 -97
rect 261 -655 266 -102
rect 1109 -577 1114 61
rect 1109 -582 1860 -577
rect 261 -660 277 -655
rect 1855 -678 1860 -582
rect 283 -683 288 -678
rect 251 -745 279 -740
rect 241 -758 275 -753
rect 231 -843 275 -838
rect 221 -856 275 -851
rect 211 -941 275 -936
rect 201 -954 275 -949
rect 191 -1039 275 -1034
rect 181 -1052 275 -1047
rect 171 -1137 275 -1132
rect 161 -1150 275 -1145
rect 151 -1235 275 -1230
rect 968 -2991 973 -1871
rect 968 -3376 973 -2996
rect 968 -3421 973 -3381
rect 977 -2924 982 -1871
rect 977 -3247 982 -2929
rect 977 -3421 982 -3252
rect 986 -2893 991 -1871
rect 986 -3118 991 -2898
rect 986 -3269 991 -3123
rect 995 -2826 1000 -1871
rect 995 -2972 1000 -2831
rect 995 -3269 1000 -2977
rect 986 -3274 1000 -3269
rect 986 -3421 991 -3274
rect 995 -3421 1000 -3274
rect 1004 -2795 1009 -1871
rect 1004 -2860 1009 -2800
rect 1004 -3421 1009 -2865
rect 1013 -2728 1018 -1871
rect 1013 -2739 1018 -2733
rect 1013 -3421 1018 -2744
rect 1022 -2602 1027 -1871
rect 1022 -2697 1027 -2607
rect 1022 -3421 1027 -2702
rect 1031 -2473 1036 -1871
rect 1031 -2630 1036 -2478
rect 1031 -3421 1036 -2635
rect 1213 -3542 1218 -2982
rect 4 -3547 1218 -3542
<< m345contact >>
rect 27 61 32 66
<< m5contact >>
rect 278 -683 283 -678
<< metal5 >>
rect 22 -678 27 66
rect 22 -683 278 -678
use stage1  stage1_0
array 0 1 1072 0 0 0
timestamp 1702538072
transform 1 0 4 0 1 1703
box 0 -1701 1068 1758
use stage2  stage2_0
timestamp 1702512363
transform 1 0 280 0 1 -1243
box 0 -623 792 1135
use stage2  stage2_1
timestamp 1702512363
transform -1 0 1868 0 1 -1243
box 0 -623 792 1135
use 12bitsub  12bitsub_0
timestamp 1702537836
transform -1 0 995 0 1 -3458
box -22 -138 976 1537
use stage2  stage2_2
timestamp 1702512363
transform 1 0 1205 0 1 -3013
box 0 -623 792 1135
<< labels >>
rlabel metal4 264 -646 264 -646 1 0
rlabel metal4 254 -646 254 -646 1 1
rlabel metal4 244 -659 244 -659 1 2
rlabel metal4 233 -663 233 -663 1 3
rlabel metal4 223 -663 223 -663 1 4
rlabel metal4 214 -663 214 -663 1 5
rlabel metal4 153 -666 153 -666 1 11
rlabel metal3 2043 -1223 2043 -1223 1 11
rlabel metal3 1178 -2646 1178 -2646 1 b11
rlabel metal3 1169 -2649 1169 -2649 1 10
rlabel metal3 1158 -2652 1158 -2652 1 9
rlabel metal3 1151 -2654 1151 -2654 1 8
rlabel metal3 1141 -2655 1141 -2655 1 7
rlabel metal3 1132 -2656 1132 -2656 1 6
rlabel metal3 1124 -2656 1124 -2656 1 5
rlabel metal3 1113 -2657 1113 -2657 1 4
rlabel metal3 1105 -2657 1105 -2657 1 3
rlabel metal3 1095 -2658 1095 -2658 1 2
rlabel metal3 1087 -2658 1087 -2658 1 1
rlabel metal3 1078 -2658 1078 -2658 1 0
rlabel metal3 1069 -2660 1069 -2660 1 0
rlabel metal3 1060 -2661 1060 -2661 1 1
rlabel metal3 1050 -2661 1050 -2661 1 2
rlabel metal3 1043 -2661 1043 -2661 1 3
rlabel metal4 1034 -2659 1034 -2659 1 4
rlabel metal4 1024 -2659 1024 -2659 1 5
rlabel metal4 1014 -2659 1014 -2659 1 6
rlabel metal4 1006 -2659 1006 -2659 1 7
rlabel metal4 996 -2658 996 -2658 1 8
rlabel metal4 989 -2658 989 -2658 1 9
rlabel metal4 980 -2657 980 -2657 1 10
rlabel metal4 970 -2658 970 -2658 1 11
<< end >>
