magic
tech scmos
timestamp 1702512363
<< metal1 >>
rect 180 588 304 596
rect 304 443 309 448
rect 180 294 304 302
rect 180 0 304 8
<< m2contact >>
rect 281 1047 286 1052
rect 281 900 286 905
rect 281 753 286 758
rect 281 606 286 611
rect 186 560 191 565
rect 186 521 191 526
rect 186 462 191 467
rect 281 459 286 464
rect 186 423 191 428
rect 186 364 191 369
rect 186 325 191 330
rect 281 312 286 317
rect 186 266 191 271
rect 186 227 191 232
rect 186 168 191 173
rect 281 165 286 170
rect 186 129 191 134
rect 186 70 191 75
rect 186 31 191 36
rect 281 18 286 23
rect 281 -129 286 -124
rect 281 -276 286 -271
rect 281 -423 286 -418
rect 281 -570 286 -565
<< metal2 >>
rect 186 1047 281 1052
rect 186 565 191 1047
rect 195 900 281 905
rect 195 526 200 900
rect 191 521 200 526
rect 204 753 281 758
rect 204 467 209 753
rect 191 462 209 467
rect 213 606 281 611
rect 213 428 218 606
rect 191 423 218 428
rect 222 459 281 464
rect 222 369 227 459
rect 191 364 227 369
rect 191 325 255 330
rect 250 317 255 325
rect 250 312 281 317
rect 191 266 259 271
rect 191 227 236 232
rect 191 168 218 173
rect 191 129 209 134
rect 191 70 200 75
rect 186 -565 191 31
rect 195 -418 200 70
rect 204 -271 209 129
rect 213 -124 218 168
rect 231 23 236 227
rect 254 170 259 266
rect 254 165 281 170
rect 231 18 281 23
rect 213 -129 281 -124
rect 204 -276 281 -271
rect 195 -423 281 -418
rect 186 -570 281 -565
<< m123contact >>
rect 165 591 170 596
rect 175 541 180 546
rect 175 491 180 496
rect 175 443 180 448
rect 304 506 309 511
rect 175 394 180 399
rect 304 359 309 364
rect 175 345 180 350
rect 175 296 180 301
rect 175 247 180 252
rect 175 198 180 203
rect 175 149 180 154
rect 175 100 180 105
rect 175 51 180 56
rect 165 0 170 5
rect 304 212 309 217
rect 304 63 309 68
<< metal3 >>
rect 165 496 170 591
rect 180 541 309 546
rect 304 511 309 541
rect 185 506 304 511
rect 165 491 175 496
rect 185 448 190 506
rect 180 443 190 448
rect 165 394 175 399
rect 165 301 170 394
rect 295 359 304 364
rect 295 350 300 359
rect 180 345 300 350
rect 165 296 175 301
rect 165 203 170 296
rect 180 247 210 252
rect 205 217 210 247
rect 205 212 304 217
rect 165 198 175 203
rect 180 149 284 154
rect 165 100 175 105
rect 165 5 170 100
rect 279 56 284 149
rect 290 63 304 68
rect 290 56 295 63
rect 180 51 295 56
use mux12  mux12_0
timestamp 1702336922
transform 1 0 14 0 1 0
box -14 0 177 596
use 12bitregout  12bitregout_0
timestamp 1702320260
transform 1 0 259 0 1 -623
box 0 0 533 1758
<< end >>
