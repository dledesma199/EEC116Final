magic
tech scmos
timestamp 1702148372
<< ntransistor >>
rect -6 -30 -4 -25
rect 11 -30 13 -25
<< ptransistor >>
rect -6 -2 -4 3
rect 11 -2 13 3
<< ndiffusion >>
rect -9 -30 -6 -25
rect -4 -30 11 -25
rect 13 -30 16 -25
<< pdiffusion >>
rect -9 -2 -6 3
rect -4 -2 1 3
rect 6 -2 11 3
rect 13 -2 16 3
<< ndcontact >>
rect -14 -30 -9 -25
rect 16 -30 21 -25
<< pdcontact >>
rect -14 -2 -9 3
rect 1 -2 6 3
rect 16 -2 21 3
<< polysilicon >>
rect -6 3 -4 6
rect 11 3 13 6
rect -6 -6 -4 -2
rect -6 -25 -4 -11
rect 11 -14 13 -2
rect 11 -25 13 -19
rect -6 -33 -4 -30
rect 11 -33 13 -30
<< polycontact >>
rect -9 -11 -4 -6
rect 8 -19 13 -14
<< metal1 >>
rect -19 7 26 12
rect -14 3 -9 7
rect 16 3 21 7
rect 1 -6 6 -2
rect -15 -11 -9 -6
rect 1 -11 23 -6
rect 2 -19 8 -14
rect 16 -25 21 -11
rect -14 -34 -9 -30
rect -19 -39 26 -34
<< end >>
