magic
tech scmos
timestamp 1702538072
<< metal1 >>
rect 423 1714 580 1722
rect 424 1652 581 1660
rect 423 1567 580 1575
rect 424 1505 581 1513
rect 423 1420 580 1428
rect 424 1358 581 1366
rect 423 1273 580 1281
rect 424 1211 581 1219
rect 423 1126 580 1134
rect 424 1064 581 1072
rect 423 979 580 987
rect 424 917 581 925
rect 423 832 580 840
rect 424 770 581 778
rect 423 685 580 693
rect 424 623 581 631
rect 423 538 580 546
rect 424 476 581 484
rect 423 391 580 399
rect 424 329 581 337
rect 423 244 580 252
rect 424 182 581 190
rect 423 97 580 105
rect 424 35 581 43
rect 1017 -84 1063 -80
rect 1022 -213 1054 -209
rect 1022 -342 1045 -338
rect 1022 -471 1036 -467
rect 1022 -600 1027 -596
rect 996 -1103 1022 -1098
rect 1017 -1112 1022 -1103
<< m2contact >>
rect 557 1670 562 1675
rect 557 1523 562 1528
rect 557 1376 562 1381
rect 557 1229 562 1234
rect 557 1082 562 1087
rect 557 935 562 940
rect 557 788 562 793
rect 557 641 562 646
rect 557 494 562 499
rect 557 347 562 352
rect 557 200 562 205
rect 557 53 562 58
rect 598 -34 603 -29
rect 598 -94 603 -89
rect 1014 -1245 1019 -1240
rect 1017 -1374 1022 -1369
<< metal2 >>
rect 429 1678 452 1683
rect 447 1675 452 1678
rect 447 1670 557 1675
rect 429 1528 434 1536
rect 429 1523 557 1528
rect 429 1381 434 1389
rect 429 1376 557 1381
rect 429 1234 434 1242
rect 429 1229 557 1234
rect 429 1087 434 1095
rect 429 1082 557 1087
rect 429 940 434 948
rect 429 935 557 940
rect 429 793 434 801
rect 429 788 557 793
rect 429 646 434 654
rect 429 641 557 646
rect 429 499 434 507
rect 429 494 557 499
rect 429 352 434 360
rect 429 347 557 352
rect 429 205 434 208
rect 429 200 557 205
rect 429 58 434 61
rect 429 53 557 58
rect 598 -89 603 -34
rect 987 -1179 991 -1178
rect 987 -1183 1018 -1179
rect 1014 -1240 1018 -1183
rect 978 -1313 1022 -1308
rect 1017 -1369 1022 -1313
rect 969 -1468 1022 -1463
rect 1017 -1498 1022 -1468
<< m3contact >>
rect 982 -1183 987 -1178
<< m123contact >>
rect 947 -62 952 -57
rect 1063 -84 1068 -79
rect 947 -191 952 -186
rect 1054 -213 1059 -208
rect 947 -320 952 -315
rect 1045 -342 1050 -337
rect 947 -449 952 -444
rect 1036 -471 1041 -466
rect 947 -578 952 -573
rect 1027 -600 1032 -595
rect 947 -707 952 -702
rect 1018 -729 1023 -724
rect 947 -836 952 -831
rect 1009 -858 1014 -853
rect 947 -965 952 -960
rect 1000 -987 1005 -982
rect 947 -1094 952 -1089
rect 991 -1103 996 -1098
rect 947 -1223 952 -1218
rect 973 -1313 978 -1308
rect 947 -1352 952 -1347
rect 964 -1468 969 -1463
rect 947 -1481 952 -1476
<< metal3 >>
rect 429 -1443 434 0
rect 429 -1701 434 -1448
rect 438 -1314 443 0
rect 438 -1701 443 -1319
rect 447 -1185 452 0
rect 447 -1701 452 -1190
rect 456 -1056 461 0
rect 456 -1701 461 -1061
rect 465 -927 470 0
rect 465 -1701 470 -932
rect 474 -798 479 0
rect 474 -1701 479 -803
rect 483 -669 488 0
rect 483 -1701 488 -674
rect 492 -540 497 0
rect 492 -1701 497 -545
rect 501 -411 506 1
rect 501 -1701 506 -416
rect 510 -282 515 0
rect 510 -1701 515 -287
rect 519 -153 524 0
rect 519 -1701 524 -158
rect 528 -24 533 0
rect 528 -1701 533 -29
rect 947 -57 952 -29
rect 947 -186 952 -158
rect 947 -315 952 -287
rect 947 -444 952 -416
rect 947 -573 952 -545
rect 947 -702 952 -674
rect 947 -831 952 -803
rect 947 -960 952 -932
rect 947 -1089 952 -1061
rect 947 -1218 952 -1190
rect 947 -1347 952 -1319
rect 947 -1476 952 -1448
rect 964 -1463 969 0
rect 964 -1701 969 -1468
rect 973 -1308 978 0
rect 973 -1701 978 -1313
rect 982 -1178 987 0
rect 982 -1701 987 -1183
rect 991 -1098 996 0
rect 991 -1701 996 -1103
rect 1000 -982 1005 0
rect 1000 -1701 1005 -987
rect 1009 -853 1014 0
rect 1009 -1701 1014 -858
rect 1018 -724 1023 0
rect 1018 -1701 1023 -729
rect 1027 -595 1032 0
rect 1027 -1701 1032 -600
rect 1036 -466 1041 0
rect 1036 -1701 1041 -471
rect 1045 -337 1050 1
rect 1045 -1701 1050 -342
rect 1054 -208 1059 0
rect 1054 -1701 1059 -213
rect 1063 -79 1068 0
rect 1063 -1701 1068 -84
<< m4contact >>
rect 429 -1448 434 -1443
rect 438 -1319 443 -1314
rect 447 -1190 452 -1185
rect 456 -1061 461 -1056
rect 465 -932 470 -927
rect 474 -803 479 -798
rect 483 -674 488 -669
rect 492 -545 497 -540
rect 501 -416 506 -411
rect 510 -287 515 -282
rect 519 -158 524 -153
rect 528 -29 533 -24
rect 947 -29 952 -24
rect 947 -158 952 -153
rect 947 -287 952 -282
rect 947 -416 952 -411
rect 947 -545 952 -540
rect 947 -674 952 -669
rect 947 -803 952 -798
rect 947 -932 952 -927
rect 947 -1061 952 -1056
rect 947 -1190 952 -1185
rect 947 -1319 952 -1314
rect 947 -1448 952 -1443
<< metal4 >>
rect 533 -29 947 -24
rect 524 -158 947 -153
rect 515 -287 947 -282
rect 506 -416 947 -411
rect 497 -545 947 -540
rect 488 -674 947 -669
rect 479 -803 947 -798
rect 470 -932 947 -927
rect 461 -1061 947 -1056
rect 452 -1190 947 -1185
rect 443 -1319 947 -1314
rect 434 -1448 947 -1443
use 12bitregout  12bitregout_0
array 0 1 535 0 0 1
timestamp 1702320260
transform 1 0 0 0 1 0
box 0 0 533 1758
use 12bitsub  12bitsub_0
timestamp 1702537836
transform -1 0 1024 0 1 -1558
box -22 -138 976 1537
<< end >>
