magic
tech scmos
timestamp 1702573332
<< metal1 >>
rect -80 7053 125 7061
rect -80 7052 -71 7053
rect -80 6914 -72 7052
rect 14 7009 47 7014
rect 33 6991 125 6999
rect -81 6906 125 6914
rect -80 6767 -72 6906
rect -7 6862 43 6867
rect 33 6844 125 6852
rect -80 6759 125 6767
rect -80 6620 -72 6759
rect -7 6715 54 6720
rect 0 6697 25 6705
rect 33 6697 125 6705
rect -81 6612 126 6620
rect -80 6473 -72 6612
rect -48 6568 20 6573
rect -51 6550 25 6558
rect 33 6550 125 6558
rect -80 6465 125 6473
rect -80 6326 -72 6465
rect -58 6421 0 6426
rect -45 6403 25 6411
rect 33 6403 125 6411
rect -80 6318 125 6326
rect -80 6179 -72 6318
rect -51 6274 55 6279
rect 20 6256 25 6264
rect 33 6256 125 6264
rect -80 6171 125 6179
rect -80 6032 -72 6171
rect -49 6127 49 6132
rect -4 6109 25 6117
rect 33 6109 125 6117
rect -80 6024 125 6032
rect -80 5885 -72 6024
rect -50 5980 42 5985
rect -39 5962 25 5970
rect 33 5962 125 5970
rect 16 5943 24 5962
rect -81 5877 125 5885
rect -80 5738 -72 5877
rect -48 5833 51 5838
rect -17 5815 25 5823
rect 33 5815 125 5823
rect -80 5730 126 5738
rect -80 5591 -72 5730
rect -55 5686 50 5691
rect 33 5668 125 5676
rect -80 5583 125 5591
rect -80 5444 -72 5583
rect -62 5539 57 5544
rect 17 5521 25 5529
rect 33 5521 125 5529
rect -80 5436 125 5444
rect -80 5310 -72 5436
rect -22 5392 41 5397
rect 33 5374 125 5382
rect -80 5302 138 5310
rect -80 5181 -72 5302
rect 64 5212 136 5220
rect -80 5173 136 5181
rect -80 5052 -72 5173
rect 32 5083 136 5091
rect -80 5044 136 5052
rect -80 4923 -72 5044
rect 18 5043 26 5044
rect -2 4954 18 4962
rect 26 4954 136 4962
rect -80 4915 136 4923
rect -80 4794 -72 4915
rect 28 4825 142 4833
rect -80 4786 138 4794
rect -80 4665 -72 4786
rect 21 4696 138 4704
rect -80 4657 136 4665
rect -80 4536 -72 4657
rect 20 4567 136 4575
rect -80 4528 136 4536
rect -80 4407 -72 4528
rect 17 4446 25 4483
rect -19 4438 136 4446
rect -80 4399 136 4407
rect -80 4278 -72 4399
rect 19 4317 27 4345
rect 5 4309 138 4317
rect -80 4270 140 4278
rect -80 4149 -72 4270
rect 17 4188 25 4207
rect -6 4180 146 4188
rect -80 4141 136 4149
rect -80 4020 -72 4141
rect 15 4059 23 4069
rect 0 4051 136 4059
rect -80 4012 136 4020
rect -80 3891 -72 4012
rect 18 3930 30 3931
rect -7 3922 136 3930
rect -80 3883 136 3891
rect -80 3753 -72 3883
rect -9 3793 18 3801
rect 26 3793 136 3801
rect -80 3745 136 3753
rect -80 3492 -72 3745
rect 26 3655 136 3663
rect -80 3484 660 3492
rect -80 3345 -72 3484
rect 156 3422 660 3430
rect -80 3337 660 3345
rect -80 3198 -72 3337
rect 74 3275 660 3283
rect -80 3190 660 3198
rect -80 3051 -72 3190
rect -40 3135 661 3136
rect -33 3128 661 3135
rect -80 3043 660 3051
rect -80 2940 -72 3043
rect 215 2981 356 2989
rect -80 2932 356 2940
rect -80 2842 -72 2932
rect 603 2896 660 2904
rect 78 2883 356 2891
rect -81 2834 356 2842
rect 596 2834 660 2842
rect -80 2744 -72 2834
rect 138 2786 140 2793
rect 148 2786 356 2793
rect 138 2785 356 2786
rect -80 2736 356 2744
rect -80 2646 -72 2736
rect 165 2688 166 2695
rect 174 2688 356 2695
rect 165 2687 356 2688
rect 596 2687 604 2834
rect 620 2749 660 2757
rect -82 2638 356 2646
rect -80 2548 -72 2638
rect 632 2602 660 2610
rect 145 2591 356 2597
rect 139 2589 356 2591
rect -80 2540 356 2548
rect 618 2540 661 2548
rect -80 2450 -72 2540
rect 621 2499 629 2540
rect 51 2491 356 2499
rect 536 2491 629 2499
rect 604 2455 670 2463
rect -80 2442 356 2450
rect -80 2316 -72 2442
rect 17 2399 356 2401
rect 23 2393 356 2399
rect -80 2308 670 2316
rect -80 2169 -72 2308
rect 61 2253 672 2254
rect 68 2246 672 2253
rect -80 2161 660 2169
rect -80 2022 -72 2161
rect 414 2099 660 2107
rect -80 2014 660 2022
rect -80 1844 -72 2014
rect 195 1952 660 1960
rect 495 1867 660 1875
rect -80 1836 259 1844
rect 495 1836 503 1867
rect -80 1707 -72 1836
rect 229 1803 248 1808
rect 598 1805 660 1813
rect 598 1766 606 1805
rect 240 1758 259 1766
rect 491 1758 606 1766
rect 2297 1722 2305 1752
rect 1962 1714 2305 1722
rect -80 1699 103 1707
rect -80 1578 -72 1699
rect 1964 1652 2086 1660
rect 26 1609 107 1617
rect -80 1570 103 1578
rect 2297 1575 2305 1714
rect -80 1449 -72 1570
rect 1963 1567 2305 1575
rect 1964 1505 2091 1513
rect 24 1480 104 1488
rect -80 1441 103 1449
rect -80 1320 -72 1441
rect 2297 1428 2305 1567
rect 1963 1420 2305 1428
rect 36 1351 107 1359
rect 1964 1358 2114 1366
rect -80 1312 108 1320
rect -80 1191 -72 1312
rect 2297 1281 2305 1420
rect 1963 1273 2305 1281
rect 5 1222 108 1230
rect 1961 1211 2088 1219
rect -80 1183 107 1191
rect -80 1062 -72 1183
rect 2297 1134 2305 1273
rect 1963 1126 2305 1134
rect -6 1093 108 1101
rect 1963 1064 2102 1072
rect -80 1054 105 1062
rect -80 933 -72 1054
rect 2297 987 2305 1126
rect 1963 979 2305 987
rect -11 964 104 972
rect -80 925 103 933
rect -80 804 -72 925
rect 1964 918 2123 925
rect 1964 917 2124 918
rect 12 835 103 843
rect 2297 840 2305 979
rect 1963 832 2305 840
rect -80 796 103 804
rect -80 675 -72 796
rect 1964 770 2128 778
rect -1 706 103 714
rect 2297 693 2305 832
rect 1963 685 2305 693
rect -80 667 103 675
rect -80 546 -72 667
rect 1963 624 2131 631
rect 1963 623 2133 624
rect -28 577 107 585
rect 2297 546 2305 685
rect -80 538 103 546
rect 1963 538 2305 546
rect -80 417 -72 538
rect 1964 476 2109 484
rect -41 448 103 456
rect -80 409 103 417
rect -80 288 -72 409
rect 2297 399 2305 538
rect 1963 391 2305 399
rect 1962 329 2124 337
rect -13 319 103 327
rect -80 280 103 288
rect -80 150 -72 280
rect 2297 252 2305 391
rect 1963 244 2305 252
rect -1 190 107 198
rect 1963 183 2129 190
rect 1963 182 2132 183
rect -80 142 109 150
rect -80 -31 -72 142
rect 2297 105 2305 244
rect 1963 97 2305 105
rect 5 52 111 60
rect 1964 35 2136 43
rect 2297 -31 2305 97
rect -80 -39 2305 -31
<< m2contact >>
rect 25 6991 33 6999
rect 25 6844 33 6852
rect 25 6697 33 6705
rect 25 6550 33 6558
rect 25 6403 33 6411
rect 25 6256 33 6264
rect 25 6109 33 6117
rect 25 5962 33 5970
rect 25 5815 33 5823
rect 25 5668 33 5676
rect 25 5521 33 5529
rect 25 5374 33 5382
rect 56 5212 64 5220
rect 24 5083 32 5091
rect 18 4954 26 4962
rect 20 4825 28 4833
rect 14 4696 21 4703
rect 12 4567 20 4576
rect 18 4483 26 4491
rect 18 4345 26 4353
rect 18 4207 26 4215
rect 18 4069 26 4077
rect 18 3931 26 3939
rect 18 3793 26 3801
rect 18 3655 26 3663
rect 148 3422 156 3430
rect 66 3275 74 3283
rect -40 3128 -33 3135
rect 207 2980 215 2989
rect 69 2883 78 2891
rect 140 2786 148 2794
rect 166 2688 174 2696
rect 139 2591 145 2597
rect 42 2491 51 2499
rect 17 2393 23 2399
rect 60 2245 68 2253
rect 406 2099 414 2107
rect 187 1952 195 1960
rect 232 1758 240 1766
rect 2086 1651 2097 1660
rect 18 1609 26 1617
rect 2091 1505 2102 1514
rect 16 1480 24 1488
rect 28 1351 36 1359
rect 2114 1357 2125 1366
rect -3 1222 5 1230
rect 2088 1212 2099 1221
rect -14 1093 -6 1101
rect 2102 1064 2113 1073
rect -19 964 -11 972
rect 2123 918 2134 927
rect 5 835 12 843
rect 2128 770 2139 779
rect -9 706 -1 714
rect 2131 624 2142 633
rect -36 577 -28 585
rect 2109 476 2120 485
rect -49 448 -41 456
rect 2124 328 2135 337
rect -21 319 -13 327
rect -9 190 -1 198
rect 2129 183 2140 192
rect -5 52 5 60
rect 2136 34 2147 43
<< metal2 >>
rect -100 6999 -92 7060
rect -100 6991 25 6999
rect -100 6852 -92 6991
rect -100 6844 25 6852
rect -100 6705 -92 6844
rect -105 6697 25 6705
rect -100 6558 -92 6697
rect -100 6550 25 6558
rect -100 6411 -92 6550
rect -103 6403 25 6411
rect -100 6264 -92 6403
rect -100 6256 25 6264
rect -100 6117 -92 6256
rect -100 6109 25 6117
rect -100 5970 -92 6109
rect -102 5962 25 5970
rect -100 5807 -92 5962
rect 17 5807 25 5823
rect -100 5799 25 5807
rect -100 5676 -92 5799
rect -100 5668 25 5676
rect -100 5529 -92 5668
rect -100 5521 25 5529
rect -100 5397 -92 5521
rect -100 5392 -72 5397
rect 1157 5392 1179 5397
rect -100 5382 -92 5392
rect 1167 5387 1172 5392
rect -100 5374 25 5382
rect -100 5220 -92 5374
rect -100 5212 56 5220
rect -100 5091 -92 5212
rect -100 5083 24 5091
rect -100 4962 -92 5083
rect -100 4954 18 4962
rect -100 4832 -92 4954
rect 13 4832 20 4833
rect -100 4825 20 4832
rect -100 4703 -92 4825
rect -100 4698 14 4703
rect -100 4574 -92 4698
rect 9 4696 14 4698
rect 5 4574 12 4576
rect -100 4567 12 4574
rect -100 4491 -92 4567
rect -100 4483 18 4491
rect -100 4353 -92 4483
rect -100 4345 18 4353
rect -100 4215 -92 4345
rect -100 4207 18 4215
rect -100 4077 -92 4207
rect -100 4069 18 4077
rect -100 3939 -92 4069
rect -100 3931 18 3939
rect -100 3801 -92 3931
rect -100 3793 18 3801
rect -100 3663 -92 3793
rect -100 3655 18 3663
rect -100 3430 -92 3655
rect 1753 3445 1758 3450
rect -100 3422 148 3430
rect -100 3283 -92 3422
rect 551 3298 556 3303
rect 1741 3298 1746 3303
rect -100 3276 66 3283
rect -100 3134 -92 3276
rect 59 3275 66 3276
rect 560 3151 565 3156
rect 1735 3151 1740 3156
rect -44 3134 -40 3135
rect -100 3130 -40 3134
rect -100 2987 -92 3130
rect -44 3128 -40 3130
rect 542 2999 547 3009
rect 569 3004 574 3009
rect 1726 3004 1731 3009
rect 200 2987 207 2989
rect -100 2980 207 2987
rect -100 2891 -92 2980
rect -100 2883 69 2891
rect -100 2793 -92 2883
rect 578 2857 583 2862
rect 1717 2857 1722 2862
rect -100 2785 140 2793
rect -100 2697 -92 2785
rect 579 2723 584 2728
rect 1700 2723 1705 2728
rect -101 2696 168 2697
rect -101 2691 166 2696
rect -100 2595 -92 2691
rect 160 2689 166 2691
rect 585 2664 590 2669
rect 1685 2664 1690 2669
rect 587 2625 592 2630
rect 1708 2625 1713 2630
rect 135 2595 139 2597
rect -100 2591 139 2595
rect -100 2497 -92 2591
rect 569 2566 574 2571
rect 1726 2566 1731 2571
rect 560 2526 565 2531
rect 1735 2527 1740 2532
rect 36 2497 42 2499
rect -100 2491 42 2497
rect -100 2398 -92 2491
rect 551 2468 556 2473
rect 1744 2468 1749 2473
rect 12 2398 17 2399
rect -100 2393 17 2398
rect -100 2253 -92 2393
rect 537 2371 542 2376
rect 1758 2368 1763 2373
rect -100 2245 60 2253
rect -100 2107 -92 2245
rect -100 2099 406 2107
rect -100 1958 -92 2099
rect 180 1958 187 1959
rect -100 1952 187 1958
rect -100 1951 188 1952
rect -100 1766 -92 1951
rect -100 1758 232 1766
rect -100 1617 -92 1758
rect 1467 1675 1472 1680
rect 2313 1660 2321 1751
rect 2097 1652 2321 1660
rect -100 1609 18 1617
rect -100 1488 -92 1609
rect 1476 1528 1481 1533
rect 2089 1505 2091 1512
rect 2313 1512 2321 1652
rect 2102 1505 2321 1512
rect 2089 1504 2321 1505
rect -100 1480 16 1488
rect -100 1359 -92 1480
rect 1485 1381 1490 1386
rect -100 1351 28 1359
rect 2313 1365 2321 1504
rect 2125 1357 2321 1365
rect -100 1230 -92 1351
rect 1494 1234 1499 1239
rect -100 1222 -3 1230
rect -100 1101 -92 1222
rect 2313 1219 2321 1357
rect 2099 1211 2321 1219
rect -100 1093 -14 1101
rect -100 971 -92 1093
rect 1504 1087 1509 1092
rect 2313 1072 2321 1211
rect 2113 1064 2321 1072
rect -26 971 -19 972
rect -100 964 -19 971
rect -100 843 -92 964
rect 1500 953 1505 958
rect 2313 926 2321 1064
rect 2134 918 2321 926
rect 1535 894 1540 899
rect 1512 855 1517 860
rect -100 836 5 843
rect -100 714 -92 836
rect -1 835 5 836
rect 1494 796 1499 801
rect 2313 779 2321 918
rect 2139 771 2321 779
rect 1485 757 1490 762
rect -100 706 -9 714
rect -100 584 -92 706
rect 1476 698 1481 703
rect 2313 633 2321 771
rect 2142 625 2321 633
rect 1462 602 1467 607
rect -41 584 -36 585
rect -101 579 -36 584
rect -100 454 -92 579
rect -41 577 -36 579
rect 2313 484 2321 625
rect 2120 476 2321 484
rect -53 454 -49 456
rect -100 450 -49 454
rect -100 324 -92 450
rect -53 448 -49 450
rect 2313 336 2321 476
rect 2135 328 2321 336
rect -26 324 -21 327
rect -100 319 -21 324
rect -100 196 -92 319
rect -15 196 -9 198
rect -100 190 -9 196
rect -100 60 -92 190
rect 1064 165 1069 233
rect 2313 190 2321 328
rect 2140 182 2321 190
rect -100 52 -5 60
rect -100 -64 -92 52
rect 2313 43 2321 182
rect 2147 35 2321 43
rect 2313 -64 2321 35
rect -100 -72 2321 -64
<< metal3 >>
rect 541 7017 546 7022
rect 1096 7017 1101 7022
rect 1625 7017 1630 7022
rect 2152 7017 2157 7022
rect 531 6870 536 6875
rect 1082 6870 1087 6875
rect 1628 6870 1633 6875
rect 2150 6870 2155 6875
rect 530 6723 535 6728
rect 1085 6723 1090 6728
rect 1615 6723 1620 6728
rect 2150 6723 2155 6728
rect 532 6576 537 6581
rect 1078 6576 1083 6581
rect 1616 6576 1621 6581
rect 2152 6576 2157 6581
rect 531 6429 536 6434
rect 1076 6429 1081 6434
rect 1614 6429 1619 6434
rect 2143 6429 2148 6434
rect 531 6282 536 6287
rect 1077 6282 1082 6287
rect 1611 6282 1616 6287
rect 2144 6282 2149 6287
rect 530 6135 535 6140
rect 1076 6135 1081 6140
rect 1611 6135 1616 6140
rect 2147 6135 2152 6140
rect 527 5988 532 5993
rect 1070 5988 1075 5993
rect 1606 5988 1611 5993
rect 2134 5988 2139 5993
rect 527 5841 532 5846
rect 1062 5841 1067 5846
rect 1598 5841 1603 5846
rect 2132 5841 2137 5846
rect 524 5694 529 5699
rect 1059 5694 1064 5699
rect 1596 5694 1601 5699
rect 2129 5694 2134 5699
rect 518 5547 523 5552
rect 1053 5547 1058 5552
rect 1590 5547 1595 5552
rect 2125 5527 2130 5532
rect 509 5384 514 5389
rect 1581 5384 1586 5389
rect 2116 5371 2121 5376
rect 1034 3643 1044 3648
rect 1969 -6 1974 0
rect 1978 -6 1983 0
rect 1987 -12 1992 0
rect 1996 -7 2001 0
rect 2005 -12 2010 0
rect 2014 -10 2019 5
rect 2023 -7 2028 0
rect 2032 -9 2037 1
rect 2041 -5 2046 0
rect 2050 -6 2055 0
rect 2059 -8 2064 0
rect 2068 -8 2073 0
<< metal4 >>
rect 1190 3690 1193 3695
rect 1294 603 1297 608
<< metal5 >>
rect 80 7106 618 7114
rect 80 7022 88 7106
rect 98 3702 103 3705
use core  core_0
timestamp 1702571561
transform 1 0 80 0 1 0
box -80 0 2140 7114
<< labels >>
rlabel metal1 -76 7057 -76 7057 1 Vdd
rlabel metal2 -95 7050 -95 7050 1 Gnd
rlabel metal1 15 7011 15 7011 1 a0
rlabel metal1 -4 6865 -4 6865 1 a1
rlabel metal1 -5 6717 -5 6717 1 a2
rlabel metal1 -46 6571 -46 6571 1 a3
rlabel metal1 -56 6424 -56 6424 1 a4
rlabel metal1 -47 6276 -47 6276 1 a5
rlabel metal1 -47 6131 -47 6131 1 a6
rlabel metal1 -44 5983 -44 5983 1 a7
rlabel metal1 -44 5836 -44 5836 1 a8
rlabel metal1 -53 5689 -53 5689 1 a9
rlabel metal1 -59 5542 -59 5542 1 aa
rlabel metal1 -20 5394 -20 5394 1 ab
rlabel metal3 1970 -4 1970 -4 1 outb
rlabel metal3 1979 -5 1979 -5 1 outa
rlabel metal3 1989 -7 1989 -7 1 out9
rlabel metal3 1997 -5 1997 -5 1 out8
rlabel metal3 2007 -8 2007 -8 1 out7
rlabel metal3 2016 -7 2016 -7 1 out6
rlabel metal3 2025 -5 2025 -5 1 out5
rlabel metal3 2034 -6 2034 -6 1 out4
rlabel metal3 2044 -2 2044 -2 1 out3
rlabel metal3 2053 -4 2053 -4 1 out2
rlabel metal3 2061 -5 2061 -5 1 out1
rlabel metal3 2070 -5 2070 -5 1 out0
rlabel metal5 100 3703 100 3703 1 sel1
rlabel metal4 1192 3691 1192 3691 1 sel2
rlabel metal4 1295 605 1295 605 1 sel3
rlabel metal2 544 3001 544 3001 1 max10
rlabel metal3 1098 7018 1098 7018 1 a20
rlabel metal3 1086 6872 1086 6872 1 a21
rlabel metal3 1086 6724 1086 6724 1 a22
rlabel metal3 1079 6578 1079 6578 1 a23
rlabel metal3 1077 6431 1077 6431 1 a24
rlabel metal3 1079 6284 1079 6284 1 a25
rlabel metal3 1078 6137 1078 6137 1 a26
rlabel metal3 1072 5990 1072 5990 1 a27
rlabel metal3 1065 5844 1065 5844 1 a28
rlabel metal3 1061 5698 1061 5698 1 a29
rlabel metal3 1054 5550 1054 5550 1 a2a
rlabel metal3 512 5385 512 5385 1 a1b
rlabel metal3 520 5551 520 5551 1 a1a
rlabel metal3 525 5695 525 5695 1 a19
rlabel metal3 528 5844 528 5844 1 a18
rlabel metal3 528 5990 528 5990 1 a17
rlabel metal3 531 6136 531 6136 1 a16
rlabel metal3 532 6286 532 6286 1 a15
rlabel metal3 533 6430 533 6430 1 a14
rlabel metal3 534 6579 534 6579 1 a13
rlabel metal3 531 6724 531 6724 1 a12
rlabel metal3 533 6873 533 6873 1 a11
rlabel metal3 542 7018 542 7018 1 a10
rlabel metal3 1627 7020 1627 7020 1 a30
rlabel metal3 1630 6872 1630 6872 1 a31
rlabel metal3 1616 6725 1616 6725 1 a32
rlabel metal3 1618 6579 1618 6579 1 a33
rlabel metal3 1616 6431 1616 6431 1 a34
rlabel metal3 1613 6285 1613 6285 1 a35
rlabel metal3 1614 6138 1614 6138 1 a36
rlabel metal3 1608 5990 1608 5990 1 a37
rlabel metal3 1600 5843 1600 5843 1 a38
rlabel metal3 1599 5696 1599 5696 1 a39
rlabel metal3 1592 5548 1592 5548 1 a3a
rlabel metal3 1582 5386 1582 5386 1 a3b
rlabel metal3 2118 5373 2118 5373 1 a4b
rlabel metal3 2129 5529 2129 5529 1 a4a
rlabel metal3 2131 5696 2131 5696 1 a49
rlabel metal3 2134 5843 2134 5843 1 a48
rlabel metal3 2136 5990 2136 5990 1 a47
rlabel metal3 2148 6137 2148 6137 1 a46
rlabel metal3 2147 6286 2147 6286 1 a45
rlabel metal3 2146 6431 2146 6431 1 a44
rlabel metal3 2155 6578 2155 6578 1 a43
rlabel metal3 2152 6725 2152 6725 1 a42
rlabel metal3 2153 6872 2153 6872 1 a41
rlabel metal3 2155 7020 2155 7020 1 a40
rlabel metal2 553 3300 553 3300 1 max11
rlabel metal2 563 3154 563 3154 1 max12
rlabel metal2 571 3008 571 3008 1 max13
rlabel metal2 579 2860 579 2860 1 max14
rlabel metal2 581 2726 581 2726 1 max15
rlabel metal2 588 2667 588 2667 1 max16
rlabel metal2 589 2627 589 2627 1 max17
rlabel metal2 571 2569 571 2569 1 max18
rlabel metal2 563 2529 563 2529 1 max19
rlabel metal2 553 2471 553 2471 1 max1a
rlabel metal2 538 2372 538 2372 1 max1b
rlabel metal2 1760 2370 1760 2370 1 max2b
rlabel metal2 1747 2471 1747 2471 1 max2a
rlabel metal2 1737 2530 1737 2530 1 max29
rlabel metal2 1728 2569 1728 2569 1 max28
rlabel metal2 1711 2628 1711 2628 1 max27
rlabel metal2 1687 2667 1687 2667 1 max26
rlabel metal2 1703 2725 1703 2725 1 max25
rlabel metal2 1719 2859 1719 2859 1 max24
rlabel metal2 1729 3006 1729 3006 1 max23
rlabel metal2 1738 3154 1738 3154 1 max22
rlabel metal2 1744 3302 1744 3302 1 max21
rlabel metal2 1755 3447 1755 3447 1 max20
rlabel metal2 1470 1678 1470 1678 1 max30
rlabel metal2 1480 1530 1480 1530 1 max31
rlabel metal2 1487 1383 1487 1383 1 max32
rlabel metal2 1497 1236 1497 1236 1 max33
rlabel metal2 1506 1089 1506 1089 1 max34
rlabel metal2 1503 956 1503 956 1 max35
rlabel metal2 1537 896 1537 896 1 max36
rlabel metal2 1514 857 1514 857 1 max37
rlabel metal2 1496 799 1496 799 1 max38
rlabel metal2 1486 760 1486 760 1 max39
rlabel metal2 1478 700 1478 700 1 max3a
rlabel metal2 1463 604 1463 604 1 max3b
rlabel metal2 1169 5389 1169 5389 1 a2b
rlabel metal1 231 1805 231 1805 1 clk
rlabel metal3 1037 3645 1037 3645 1 a2b
<< end >>
